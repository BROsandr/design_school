module simple_add_sub (
  input  [7:0] operandA, operandB,        // два входных 8-ми битных операнда
  output [15:0] out_mul, out_div, out_rem // Для умножения, чтобы избежать переполения выходная
                                          //   разрядность должна быть не меньше, чем сумма
                                          //   разрядностей операндов для беззнаковго случая и сумма
                                          //   разрядностей операндов -1 для знакового. Для данного 
                                          //   случая это 16 бит и 15 бит. Для знакового случая
                                          //   разрядность меньше из-за наличия старшего бита знака.
);
  assign out_mul = operandA * operandB; // Умножение 8 * 8 = 64
  assign out_div = operandA / operandB; // Деление 16 / 3 = 5. Округление до целого числа вниз.
  assign out_rem = operandA % operandB; // Остаток от деления 16 % 3 = 1
  // ВАЖНО. Использование операций деления и остаток от деления не используется в синтезируемом
  //   коде, только для симуляции. Так как дает очень сложную реализацию по площади и очень плохие
  //   тайминги. Например в процессорах деление реализуется итерационными алгоритмами.
endmodule
