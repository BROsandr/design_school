module simple_add_sub (
  input  [7:0] operandA, operandB, // два входных 8-ми битных операнда
  output [8:0] out_sum, out_dif    // Выходы для арифметических операций имеют дополнительный 9-й
                                   //   бит переполнения
);
  // Максимальное 8-ми битное беззнаковое число 255.
  //   При сложении 255 + 255 получится 510, которое можно представить минимум 9-ю битами.
  assign out_sum = operandA + operandB;
  assign out_dif = operandA - operandB;
  // Если сделать выход сумматора 8-ми битным, то случится переполнение и результат сложения 255 + 3
  //   будет равен 2.
endmodule
