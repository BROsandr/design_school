module top (
  input        clk,
  input  [8:0] a,
  input        b,
  output [3:0] q
);
// reg используют при поведенческом(behavioral) описании схемы.о Если регистру постоянно 
//   присваивается значение комбинаторной(логической) функции, то он ведет себя точно как провод
//   (wire). Если же регистру присваивается значение в синхронной логике, например по фронту сигнала
//   тактовой частоты, то ему, в конечном счете, будет соответствовать физический D-триггер или
//   группа D-триггеров. D-триггер - это лолгический элемент способный запоминать один бит
//   информации.
  reg [3:0] c;
endmodule
