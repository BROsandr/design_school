wire [10:0] a = 7;              // 32-х битное десятичное число, которое будет "обрезано"
wire [10:0] b = 'd7;            // 11-ти битное десятичное число
wire [10:0] b = 11'd7;          // 11-ти битное десятичное число
wire [3:0]  c = 4'b0101;        // 4-ч ибтное двоичное число
wire [3:0]  d = 8'h7B;          // 8-ми битное шестнадцатеричное число 7B
wire [47:0] e = 48'hEFCA7ED98F; // 48-ми битное шестнадцатиричное число

wire signed [10:0] b = -11'd7;  // 11-ти битное отрицательное десятичное число
