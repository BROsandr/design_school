module top (
  input            clk,
  input      [8:0] a,
  input            b,
  output reg [3:0] q // выходные сигналы и шины можно объявлять как reg
);
endmodule
